
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
use std.textio.all;
use work.txt_util.all;

ENTITY testbench IS
END testbench;
 
ARCHITECTURE behavior OF testbench IS
 
  --Inputs
  signal CLK : std_logic := '0';
  signal RST : std_logic := '0';
  signal START : std_logic := '0';
  signal PLAIN : std_logic_vector(127 downto 0) := (others => '0');
  signal KEY : std_logic_vector(127 downto 0) := (others => '0');

  --Outputs
  signal CIPHER : std_logic_vector(127 downto 0);
  signal DONE : std_logic;

  -- Clock period definitions
  constant CLK_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   AES_INST: entity work.AES_128_ENC PORT MAP (
          CLK => CLK,
          RST => RST,
          START => START,
          PLAIN => PLAIN,
          KEY => KEY,
          CIPHER => CIPHER,
          DONE => DONE
        );

   -- Clock process definitions
   CLK_process :process
   begin
		CLK <= '0';
		wait for CLK_period/2;
		CLK <= '1';
		wait for CLK_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
    type test_cases_type is array(0 to 256) of std_logic_vector(127 downto 0);
    constant test_cleartexts : test_cases_type := (
      (x"32" & x"43" & x"f6" & x"a8" & x"88" & x"5a" & x"30" & x"8d" & x"31" & x"31" & x"98" & x"a2" & x"e0" & x"37" & x"07" & x"34"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00")
      );
    constant test_keys : test_cases_type := (
      (x"2b" & x"7e" & x"15" & x"16" & x"28" & x"ae" & x"d2" & x"a6" & x"ab" & x"f7" & x"15" & x"88" & x"09" & x"cf" & x"4f" & x"3c"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"01"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"03"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"07"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"0f"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"1f"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"3f"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"7f"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"01" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"03" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"07" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"0f" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"1f" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"3f" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"7f" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"01" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"03" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"07" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"0f" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"1f" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"3f" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"7f" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"01" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"03" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"07" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"0f" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"1f" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"3f" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"7f" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"01" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"03" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"07" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"0f" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"1f" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"3f" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"7f" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"01" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"03" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"07" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"0f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"1f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"3f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"7f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"01" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"03" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"07" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"0f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"1f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"3f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"7f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"01" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"03" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"07" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"0f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"1f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"3f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"7f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"01" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"03" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"07" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"0f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"1f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"3f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"7f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"01" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"03" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"07" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"0f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"1f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"3f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"7f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"01" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"03" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"07" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"0f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"1f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"3f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"7f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"00" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"01" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"03" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"07" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"0f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"1f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"3f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"7f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"00" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"01" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"03" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"07" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"0f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"1f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"3f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"7f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"00" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"01" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"03" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"07" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"0f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"1f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"3f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"7f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"00" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"01" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"03" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"07" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"0f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"1f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"3f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"7f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"00" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"01" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"03" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"07" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"0f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"1f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"3f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"7f" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fe"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fc"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f8"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f0"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"e0"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"c0"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"80"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fe" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fc" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f8" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f0" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"e0" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"c0" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"80" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fe" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fc" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f8" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f0" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"e0" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"c0" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"80" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fe" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fc" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f8" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f0" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"e0" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"c0" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"80" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fe" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fc" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f8" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f0" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"e0" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"c0" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"80" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fe" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fc" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f8" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f0" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"e0" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"c0" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"80" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fe" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fc" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f8" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"e0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"c0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"80" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fe" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fc" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f8" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"e0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"c0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"80" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fe" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fc" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f8" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"e0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"c0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"80" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fe" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fc" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f8" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"e0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"c0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"80" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fe" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"fc" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f8" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"f0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"e0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"c0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"80" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"ff" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"fe" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"fc" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"f8" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"f0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"e0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"c0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"80" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"ff" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"fe" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"fc" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"f8" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"f0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"e0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"c0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"80" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"ff" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"fe" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"fc" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"f8" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"f0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"e0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"c0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"80" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"ff" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"fe" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"fc" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"f8" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"f0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"e0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"c0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"80" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"ff" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"fe" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"fc" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"f8" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"f0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"e0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"c0" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00"),
      (x"80" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00" & x"00")
      );
    variable l: line;
    file log_file : text;
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
      RST <= '1';
      wait for CLK_period*10;
      RST <= '0';
      
      -- insert stimulus here
      --file_open(log_file,"D:\testbench.log",write_mode);
      for i in 0 to 256 loop
        KEY <= test_keys(i);
        PLAIN <= test_cleartexts(i);
        wait for CLK_period*2;
        START <= '1';
        wait for CLK_period*2;
        START <= '0';
        wait until DONE = '1';
        report hstr(CIPHER);
        --write(l, to_lower(hstr(CIPHER)));
        --writeline(log_file, l);
        wait for CLK_period*2;
      end loop;
      --file_close(log_file);
      
      wait;
   end process;

END;
